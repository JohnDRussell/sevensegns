-----------------------------------------
---- SevenSegNS_tb.vhdl
---- Seven segment driver with 4 input
---- buttons

---- Author: Derby Russell
---- Date: 12-13-2013
-----------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.ALL;

entity sevensegns_tb is
end sevensegns_tb;

architecture behavioral_3 of sevensegns_tb is
    component main_7_seg
     port(b1,b2,b3,b4 : in std_logic;
          clk         : in std_logic;
          sseg        : out std_logic_vector(0 to 6);
          anodes      : out std_logic_vector (3 downto 0);
          reset       : in std_logic
          );
    end component;
    for sevensegns_0: main_7_seg use entity work.main_7_seg;
    signal b1 : std_logic; 
    signal b2 : std_logic; 
    signal b3 : std_logic; 
    signal b4 : std_logic; 
    signal clk : std_logic; 
    signal sseg : std_logic_vector (0 to 6); 
    signal anodes : std_logic_vector (3 downto 0); 
    signal reset : std_logic;
begin
    -- Component instantiation.
    sevensegns_0: main_7_seg port map (b1 => b1, b2 => b2, b3 => b3,
                                       b4 => b4, clk => clk,
                                       sseg => sseg, anodes => anodes,
                                       reset => reset);

    process
        type pattern_type is record
        -- The inputs of the main_7_seg.
        b1a, b2a, b3a, b4a, clka, reseta : std_logic;
        -- The expected outputs of the main_7_seg.
        -- sseg, anodes : std_logic_vector (0 to 6) ;
        -- anodes : std_logic_vector (3 to 0);
        end record;
        -- The patterns to apply.
        type pattern_array is array (natural range <>) of pattern_type;
        constant patterns : pattern_array :=
          (('0', '0', '0', '0', '1', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '1', '1'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('1', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('1', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('1', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('1', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('1', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('1', '0', '0', '0', '0', '0'), -- button 1 is done
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '1', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '1', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '1', '0', '0', '0'),
           ('0', '0', '1', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '1', '0', '0'),
           ('0', '0', '0', '1', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '0'),
           ('0', '0', '0', '0', '1', '0'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '1', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'),
           ('0', '0', '0', '0', '0', '1'));
    begin
       -- Check each pattern.
       for i in patterns'range loop
          -- Set the inputs.
          b1 <= patterns(i).b1a;
          b2 <= patterns(i).b2a;
          b3 <= patterns(i).b3a;
          b4 <= patterns(i).b4a;
          clk <= patterns(i).clka;
          reset <= patterns(i).reseta;
          -- Wait for the results.
          wait for 1 ns;
          -- Check the outputs.
          if sseg = "0000001" then
              report "sseg value 0000001" severity error;
          elsif sseg = "1001111" then
              report "sseg value 1001111" severity error;
          elsif sseg = "0010010" then
              report "sseg value 0010010" severity error;
          elsif sseg = "0000110" then
              report "sseg value 0000110" severity error;
          elsif sseg = "1001100" then
              report "sseg value 1001100" severity error;
          elsif sseg = "0100100" then
              report "sseg value 0100100" severity error;
          elsif sseg = "0100000" then
              report "sseg value 0100000" severity error;
          elsif sseg = "0001111" then
              report "sseg value 0001111" severity error;
          elsif sseg = "0000000" then
              report "sseg value 0000000" severity error;
          elsif sseg = "0000100" then
              report "sseg value 0000100" severity error;
          else
              report "sseg value 0010000" severity error;
          end if;

          if anodes = "1110" then
              report "anodes value 1110" severity error;
          elsif anodes = "1101" then
              report "anodes value 1101" severity error;
          elsif anodes = "1011" then
              report "anodes value 1011" severity error;
          elsif anodes = "0111" then
              report "anodes value 0111" severity error;
          else
              report "anodes value null" severity error;
          end if;
       end loop;
       assert false report "end of test" severity note;
       -- Wait forever; this will finish the simulation.
       wait;
    end process;
end behavioral_3;




